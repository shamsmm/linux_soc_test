module gpio_wrapped(slave_bus_if.slave bus)

endmodule